module main
fn main(){
	f0()
	f1()
	f2()
}
