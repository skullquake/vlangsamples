module d
pub fn f2(){
	println('f2:start')
	println('f2:end')
}
