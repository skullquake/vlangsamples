module main
import c
import d
fn main(){
	f0()
	c.f1()
	d.f2()
}
