module c
pub fn f1(){
	println('f1:start')
	println('f1:end')
}
